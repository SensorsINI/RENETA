
import definesPkg::*;

// SMEM Read Request Generator (CH_S0)
//   For fetching NZI

// cfg_ready initialized to 1?
//           set to 1 only when cfg_valid==1?

// Modified for dtv1.0_perf_estm:
//   Set ready_i_nzn=0 when pop_nzn if empty
//     Set rd_avalid to 0 when waiting for ready_i_nzn after a completed read address transaction
//   PROC_MTxV_SP: send request for reading NZI for cnt1 == 0 to cfg_cnt1_r,
//     for simpler IPM_DRG pop_nzi logic.
//     Should set cfg_cnt1_r = 0 in the future to avoid sending redundant requests.


module IPM_SRG0 #(
    // parameter NUM_PE        = 16,               //16
    // parameter MAX_N         = 256,              //1024
    // parameter MAX_M         = 256,              //32
    // parameter MAX_NoP       = MAX_N/NUM_PE,     //64

    parameter SMEM_WW       = 16,
    parameter SMEM_DEPTH    = MAX_M*MAX_NoP*4,

    localparam ADDR_BW      = $clog2(SMEM_DEPTH),       // MSB: bank(SRAM0/SRAM1)
    localparam WSEL_BW      = $clog2(NUM_PE) + 1        // {WordOp, WordIdx}
    // localparam NZL_HA_BW    = $clog2(MAX_NoP*MAX_M),    // NZL head address bit-width
    // localparam MAX_CNT      = (MAX_N>MAX_M)? (MAX_N):(MAX_M)
) (
    input  logic                        clk,
    input  logic                        rstn,
    
    input  logic                        cfg_valid,
    // input  PROC_t                       cfg_proc,
    // input  logic [$clog2(MAX_CNT)-1:0]  cfg_cnt0,
    // input  logic [$clog2(MAX_CNT)-1:0]  cfg_cnt1,
    // input  logic [$clog2(MAX_CNT)-1:0]  cfg_cnt2,
    input  cfg_t                        cfg_data,
    output logic                        cfg_ready,

    input  logic [ADDR_BW-1:0]          smem_addr0,
    input  logic [NZL_HA_BW-1:0]        nzl_head_addr,
    input  logic [$clog2(NUM_PE)-1:0]   nzl_head_peid,

    input  logic [$clog2(MAX_N)-1:0]    din_nzn,
    output logic                        pop_nzn,
    input  logic                        empty_nzn,

    // ---------------- SMEM Read Channels ----------------
    output logic [WSEL_BW-1:0]          rd_wsel   [0:0],
    output logic [ADDR_BW-1:0]          rd_addr   [0:0],
    output logic                        rd_avalid [0:0],
    input  logic                        rd_aready [0:0]
    // input  logic [SMEM_WW-1:0]          rd_dout   [0:0][0:NUM_PE-1],
    // input  logic                        rd_dvalid [0:0][0:NUM_PE-1],
    // output logic                        rd_dready [0:0]
    
);


// -----------------------------------------------------------------------------
// Global variables

    // Overall - control signals
    logic                               rstn_init;
    
    // Overall - flags
    logic [0:1]                         f_O;
    logic [0:1]                         f_O_rd0;
    
    // Input Signal
    PROC_t                              cfg_proc_r;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt0_r;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt1_r;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt2_r;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt0_r1;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt1_r1;
    logic [$clog2(MAX_CNT)-1:0]         cfg_cnt2_r1;

    logic [ADDR_BW-1:0]                 smem_addr0_r;
    logic [NZL_HA_BW-1:0]               nzl_head_addr_r;
    logic [$clog2(NUM_PE)-1:0]          nzl_head_peid_r;

    // logic [$clog2(MAX_N)-1:0]           din_nzn_r;
    // logic [0:1]                         pop_nzn_r;

    logic                               ready_i_eff;
    logic                               ready_i_nzn;

    // Output Signal
    logic [0:1]                         valid_o_r;
    logic [WSEL_BW-1:0]                 rd_wsel_r   [0:0];
    logic [ADDR_BW-1:0]                 rd_addr_r   [0:0];
    logic                               rd_avalid_r0[0:0];
    logic                               rd_avalid_r1[0:0];
    logic                               rd_aready_d [0:0];
    
    // FSM - states
    // (* mark_debug = "true" *)
    enum logic [1:0] {S_IDLE, S_INIT, S_GEN} state;
    logic                               f_proc_end;
    
    // SMEM Data I/O Counters
    logic [$clog2(MAX_CNT)-1:0]         cnt0;   // Inner most loop
    logic [$clog2(MAX_CNT)-1:0]         cnt1;
    logic [$clog2(MAX_CNT)-1:0]         cnt2;   // Outer most loop
    logic                               f_cnt_o;
    logic [0:1]                         f_cnt_o_r;

    // NZL Address Counters
    logic [NZL_HA_BW-1:0]               nzi_addr;       // MxV_SP, VXV_SP
    logic [$clog2(NUM_PE)-1:0]          nzi_peid;
    logic [NZL_HA_BW-1:0]               nzi_addr2;      // MTxV_SP
    logic [$clog2(NUM_PE)-1:0]          nzi_peid2;
    
    
// -----------------------------------------------------------------------------
// Module body

    
    // FSM
    always_ff @(posedge clk) begin
        if (!rstn) begin
            state <= S_IDLE;
        end else begin
            case (state) inside
    
                S_IDLE : begin              // Idle
                    if (cfg_valid) begin
                        state <= S_INIT;
                    end
                end
                
                S_INIT : begin              // Initialize
                    if (cfg_proc_r inside {PROC_MxV_SP, PROC_MTxV_SP, PROC_VXV_SP})
                        state <= S_GEN;
                    else
                        state <= S_IDLE;
                end
                
                S_GEN : begin
                    if (f_proc_end) begin
                        state <= S_IDLE;
                    end
                end

                default : begin
                    state <= S_IDLE;
                end

            endcase
        end
    end

    assign f_proc_end = f_cnt_o_r[1] && valid_o_r[1] && ready_i_eff;
    
    
    
    // Configure Signals

    always_ff @(posedge clk) begin
        if (!rstn) begin
            cfg_ready <= 1'b1;
        end else begin
            case (state) inside
                // // Assert when there is a valid cfg. Deassert at the next cc.
                // // Should be initialized to 0.
                // S_IDLE : begin
                //     if (cfg_valid) begin
                //         cfg_ready <= 1'b1;
                //     end
                // end
                // ???: Deassert when a procedure is started
                S_IDLE : begin
                    if (cfg_valid) begin
                        cfg_ready <= 1'b0;
                    end
                end
                // Assert when a procedure is finished
                S_GEN : begin
                    if (f_proc_end) begin
                        cfg_ready <= 1'b1;
                    end
                end
                default : begin
                    cfg_ready <= 1'b0;
                end
            endcase
        end
    end

    always_ff @(posedge clk) begin
        if (!rstn) begin
            cfg_proc_r <= PROC_IDLE;
        end else begin
            case (state) inside
                S_IDLE : begin
                    if (cfg_valid) begin
                        cfg_proc_r <= cfg_data.proc;
                    end
                end
                S_INIT : begin
                    if (!(cfg_proc_r inside {PROC_MxV_SP, PROC_MTxV_SP, PROC_VXV_SP})) begin
                        cfg_proc_r <= PROC_IDLE;
                    end
                end
                S_GEN : begin
                    if (f_proc_end) begin
                        cfg_proc_r <= PROC_IDLE;
                    end
                end
                default : begin
                    cfg_proc_r <= cfg_proc_r;
                end
            endcase
        end
    end

    always_ff @(posedge clk) begin
        if (!rstn) begin
            cfg_cnt0_r1     <= '0;
            cfg_cnt1_r1     <= '0;
            cfg_cnt2_r1     <= '0;
            smem_addr0_r    <= '0;
            nzl_head_addr_r <= '0;
            nzl_head_peid_r <= '0;
        end else if ((state == S_IDLE) && cfg_valid) begin
            cfg_cnt0_r1     <= cfg_data.cnt0;
            cfg_cnt1_r1     <= cfg_data.cnt1;
            cfg_cnt2_r1     <= cfg_data.cnt2;
            smem_addr0_r    <= smem_addr0;
            nzl_head_addr_r <= nzl_head_addr;
            nzl_head_peid_r <= nzl_head_peid;
        end
    end

    always_ff @(posedge clk) begin
        if (!rstn) begin
            cfg_cnt0_r <= '0;
            cfg_cnt1_r <= '0;
            cfg_cnt2_r <= '0;
        end else begin
            case (cfg_proc_r) inside
                PROC_MxV_SP : begin
                    if (state == S_INIT) begin
                        cfg_cnt0_r <= cfg_cnt0_r1;
                        cfg_cnt1_r <= din_nzn;
                        cfg_cnt2_r <= cfg_cnt2_r1;
                    end
                end
                PROC_MTxV_SP : begin
                    if (state == S_INIT) begin
                        cfg_cnt0_r <= cfg_cnt0_r1;
                        cfg_cnt1_r <= cfg_cnt1_r1;
                        cfg_cnt2_r <= din_nzn;
                    end
                end
                PROC_VXV_SP : begin
                    if (state == S_INIT) begin
                        cfg_cnt0_r <= din_nzn;
                        cfg_cnt1_r <= cfg_cnt1_r1;
                        cfg_cnt2_r <= cfg_cnt2_r1;
                    end else if (valid_o_r[0] && (cnt0 == cfg_cnt0_r) && !f_cnt_o && ready_i_eff) begin
                        cfg_cnt0_r <= din_nzn;
                    end
                end
                default : begin
                    if (state == S_INIT) begin
                        cfg_cnt0_r <= cfg_cnt0_r1;
                        cfg_cnt1_r <= cfg_cnt1_r1;
                        cfg_cnt2_r <= cfg_cnt2_r1;
                    end
                end
            endcase
        end
    end

    // (!) Not registered
    // (!) No empty check
    always_comb begin
        pop_nzn = 1'b0;
        case (cfg_proc_r) inside
            PROC_MxV_SP : begin
                if (state == S_INIT) begin
                    pop_nzn = 1'b1;
                end
            end
            PROC_MTxV_SP : begin
                if (state == S_INIT) begin
                    pop_nzn = 1'b1;
                end
            end
            PROC_VXV_SP : begin
                if (state == S_INIT) begin
                    pop_nzn = 1'b1;
                end else if (valid_o_r[0] && (cnt0 == cfg_cnt0_r) && !f_cnt_o && ready_i_eff) begin   // S_GEN
                    pop_nzn = 1'b1;
                end
            end
            default : begin
                if (state == S_INIT) begin
                    pop_nzn = 1'b0;
                end
            end
        endcase
    end



    // Control Signals
    
    // assign ready_i_eff = rd_aready[0];  // TODO
    assign ready_i_eff = rd_aready[0] && ready_i_nzn;

    always_comb begin
        case (cfg_proc_r) inside
            PROC_MxV_SP, PROC_MTxV_SP : begin
                ready_i_nzn = 1'b1;
            end
            PROC_VXV_SP : begin
                ready_i_nzn = 1'b1;
                if (valid_o_r[0] && (cnt0 == cfg_cnt0_r) && !f_cnt_o && empty_nzn)
                    ready_i_nzn = 1'b0;
            end
            default : begin 
                ready_i_nzn = 1'b1;
            end
        endcase
    end

    assign valid_o_r[0] = f_O[0];
    always_ff @(posedge clk) begin
        if (!rstn || !rstn_init) begin
            valid_o_r[1] <= 1'b0;
        end else if (ready_i_eff) begin
            valid_o_r[1] <= valid_o_r[0];
        end
    end
    


    // assign rstn_init = !(state == S_INIT);
    always_ff @(posedge clk) begin
        if (!rstn) begin
            rstn_init <= 1'b1;
        end else begin
            if ((state == S_IDLE) && cfg_valid) begin
                rstn_init <= 1'b0;
            end else begin
                rstn_init <= 1'b1;
            end
        end
    end
    
    
    
    // Flags

    // Flag - Overall output
    always_ff @(posedge clk) begin
        if (!rstn) begin
            f_O[0] <= 1'b0;
        end else begin
            case (state) inside
                // Assert at transition S_INIT -> S_GEN
                S_INIT : begin
                    if (cfg_proc_r inside {PROC_MxV_SP, PROC_MTxV_SP, PROC_VXV_SP}) begin
                        f_O[0] <= 1'b1;
                    end
                end
                // Deassert at transition S_GEN -> S_IDLE
                S_GEN : begin
                    if (f_cnt_o_r[0] && valid_o_r[0] && ready_i_eff) begin
                        f_O[0] <= 1'b0;
                    end
                end
                default : begin
                    f_O[0] <= 1'b0;
                end
            endcase
        end
    end
    
    always_ff @(posedge clk) begin
        if (!rstn || !rstn_init) begin
            f_O[1] <= '0;
        end else if ((valid_o_r[0] || valid_o_r[1]) && ready_i_eff) begin
            f_O[1] <= f_O[0];
        end
    end
    
    // Flag - SMEM Read Channel 1
    always_ff @(posedge clk) begin
        if (!rstn) begin
            f_O_rd0[0] <= 1'b0;
        end else begin
            case (state) inside
                // Assert at transition S_INIT -> S_GEN
                S_INIT : begin
                    case (cfg_proc_r) inside
                        PROC_MxV_SP, PROC_MTxV_SP, PROC_VXV_SP : f_O_rd0[0] <= 1'b1;
                        default                                : f_O_rd0[0] <= 1'b0;
                    endcase
                end
                // Deassert at transition S_GEN -> S_IDLE
                S_GEN : begin
                    if (f_cnt_o_r[0] && valid_o_r[0] && ready_i_eff) begin
                        f_O_rd0[0] <= 1'b0;
                    end
                end
                default : begin
                    f_O_rd0[0] <= 1'b0;
                end
            endcase
        end
    end
    
    always_ff @(posedge clk) begin
        if (!rstn || !rstn_init) begin
            f_O_rd0[1] <= '0;
        end else if ((valid_o_r[0] || valid_o_r[1]) && ready_i_eff) begin
            f_O_rd0[1] <= f_O_rd0[0];
        end
    end
    
    
    
    // SMEM Data Counters
    always_ff @(posedge clk) begin
        if (!rstn || !rstn_init) begin
            cnt0 <= 0;
            cnt1 <= 0;
            cnt2 <= 0;
        end else if (valid_o_r[0] && ready_i_eff) begin
            if (cnt0 == cfg_cnt0_r) begin
                if (cnt1 == cfg_cnt1_r) begin
                    if (cnt2 == cfg_cnt2_r) begin
                        cnt2 <= 0;
                    end else begin
                        cnt2 <= cnt2 + 1;
                    end
                    cnt1 <= 0;
                end else begin
                    cnt1 <= cnt1 + 1;
                end
                cnt0 <= 0;
            end else begin
                cnt0 <= cnt0 + 1;
            end
        end
    end
    
    assign f_cnt_o = (cnt2 == cfg_cnt2_r) && (cnt1 == cfg_cnt1_r) && (cnt0 == cfg_cnt0_r);
    
    assign f_cnt_o_r[0] = f_cnt_o && valid_o_r[0];
    always_ff @(posedge clk) begin
        if (!rstn || !rstn_init) begin
            f_cnt_o_r[1] <= '0;
        end else if ((valid_o_r[0] || valid_o_r[1]) && ready_i_eff) begin
            f_cnt_o_r[1] <= f_cnt_o_r[0];
        end
    end
    
    
    // NZL address counters
    always_ff @(posedge clk) begin
        // if (!rstn) begin
        //     nzi_addr <= '0;
        //     nzi_peid <= '0;
        // end else
        if (!rstn_init) begin
            nzi_addr <= nzl_head_addr_r;
            nzi_peid <= nzl_head_peid_r;
        end else if (valid_o_r[0] && ready_i_eff) begin     // MxV_SP, VXV_SP
            if ((cnt1 == cfg_cnt1_r) && (cnt0 == cfg_cnt0_r)) begin
                nzi_addr <= nzl_head_addr_r;
                nzi_peid <= nzl_head_peid_r;
            end else begin
                if (nzi_peid == '1) begin
                    nzi_addr <= nzi_addr + 1;
                end
                nzi_peid <= nzi_peid + 1;
            end
        end
    end
    
    always_ff @(posedge clk) begin
        // if (!rstn) begin
        //     nzi_addr2 <= '0;
        //     nzi_peid2 <= '0;
        // end else
        if (!rstn_init) begin
            nzi_addr2 <= nzl_head_addr_r;
            nzi_peid2 <= nzl_head_peid_r;
        // end else if (valid_o_r[0] && (cnt1 == 0) && ready_i_eff) begin     // MTxV_SP
        end else if (valid_o_r[0] && (cnt1 == cfg_cnt1_r) && ready_i_eff) begin // MTxV_SP
            // && (cnt0 == 0)
            if (nzi_peid2 == '1) begin
                nzi_addr2 <= nzi_addr2 + 1;
            end
            nzi_peid2 <= nzi_peid2 + 1;
        end
    end
    


    // SMEM Read Channel 0 - read request signals
    always_comb begin
        case (cfg_proc_r)
            PROC_MxV_SP : begin
                rd_avalid_r0[0] = f_O_rd0[0];
                rd_wsel_r[0] = {1'b1, nzi_peid};
                rd_addr_r[0] = smem_addr0_r + nzi_addr;
            end
            PROC_MTxV_SP : begin
                rd_avalid_r0[0] = f_O_rd0[0]; // && (cnt1 == 0);
                rd_wsel_r[0] = {1'b1, nzi_peid2};
                rd_addr_r[0] = smem_addr0_r + nzi_addr2;
            end
            PROC_VXV_SP : begin
                rd_avalid_r0[0] = f_O_rd0[0];
                rd_wsel_r[0] = {1'b1, nzi_peid};
                rd_addr_r[0] = smem_addr0_r + nzi_addr;
            end

            default : begin
                rd_avalid_r0[0] = 1'b0;
                rd_wsel_r[0] = '0;
                rd_addr_r[0] = '0;
            end
        endcase
    end
    
    always_ff @(posedge clk) begin
        for (int unsigned ch_idx = 0; ch_idx <= 0; ch_idx++) begin
            if (!rstn || !rstn_init) begin
                rd_avalid_r1[ch_idx] <= '0;
                rd_wsel[ch_idx] <= '0;
                rd_addr[ch_idx] <= '0;
            end else if (ready_i_eff) begin
                rd_avalid_r1[ch_idx] <= rd_avalid_r0[ch_idx];
                if (rd_avalid_r0[ch_idx]) begin
                    rd_wsel[ch_idx] <= rd_wsel_r[ch_idx];
                    rd_addr[ch_idx] <= rd_addr_r[ch_idx];
                end
            end
        end
    end

    // Set rd_avalid to 0 when waiting for ready_i_nzn after a completed read address transaction
    always_ff @(posedge clk) begin
        if (!rstn) begin
            rd_aready_d[0] <= 1'b0;
        end else begin
            if (ready_i_eff) begin
                rd_aready_d[0] <= 1'b0;
            end else begin
                rd_aready_d[0] <= rd_aready_d[0] || (rd_avalid[0] && rd_aready[0]);
            end
        end
    end

    assign rd_avalid[0] = rd_avalid_r1[0] && !rd_aready_d[0];



endmodule
